library verilog;
use verilog.vl_types.all;
entity Generator_vlg_vec_tst is
end Generator_vlg_vec_tst;
